library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Intro is

	port 
	(
		a	   : in std_logic;
		b	   : in std_logic;
		result : out std_logic
	);

end entity;

architecture rtl of Intro is
begin

	result <= a and b;

end rtl;
